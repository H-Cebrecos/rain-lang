entity uart_rx is
generic
(
	G_DATA_BITS	: natural := 8,
	G_PARITY	: parity_none,
	G_STOP_BITS	: natural_range_1_to_2
);
port
(
	clk	: In  std_logic,
	rst	: In  std_logic,
	rx	: In  std_logic,
	data	: Out std_logic_vector(7 downto 0),
	valid	: Out std_logic,
	frame_err	: Out std_logic,
	parity_err	: Out std_logic
);
end uart_rx;

architecture implementation of uart_rx is
	-- declarations
begin
	-- contents
-- Autogenerated asynchronously asserted, synchronously deasserted signal synchronizer.
process ({clk}, rst)
begin
    if rst = '1' then
        sync1_sync_stages <= (others => '1');
    elsif rising_edge({{clk}}) then
        sync1_sync_stages(1) <= '0';
        for i in 2 to sync1_STAGES loop
            sync1_sync_stages(i) <= sync1_sync_stages(i-1);
        end loop;
    end if;
end process;

rst_out <= sync1_sync_stages(sync1_STAGES)

-- ASYNC_REG attribute on each flip-flop
for i in 1 to sync1_STAGES generate
    attribute ASYNC_REG : string;
    attribute ASYNC_REG of sync1_sync_stages(i) : signal is "TRUE";
end generate;
-- End of Sync-Async synchronizer.
end implementation;

